** Profile: "SCHEMATIC1-021"  [ e:\�q�u���\1______________________�@�~\chapther2\021\p021\021-schematic1-021.sim ] 

** Creating circuit file "021-schematic1-021.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\pwrmos.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 101 0.1 10e8
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\021-SCHEMATIC1.net" 


.END
