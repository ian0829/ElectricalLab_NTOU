** Profile: "SCHEMATIC1-test"  [ C:\1________________________\CHAPTHER2\021\test\test-SCHEMATIC1-test.sim ] 

** Creating circuit file "test-SCHEMATIC1-test.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1m 0 50n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\test-SCHEMATIC1.net" 


.END
