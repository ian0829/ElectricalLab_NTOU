** Profile: "SCHEMATIC1-092_2"  [ C:\1________________________\chapther2\091\091_2-schematic1-092_2.sim ] 

** Creating circuit file "091_2-schematic1-092_2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\siemens.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 101 0.1 10e9
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\091_2-SCHEMATIC1.net" 


.END
