** Profile: "SCHEMATIC1-051"  [ C:\1________________________\chapther2\051\051-SCHEMATIC1-051.sim ] 

** Creating circuit file "051-SCHEMATIC1-051.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.5m 0 50n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\051-SCHEMATIC1.net" 


.END
