** Profile: "SCHEMATIC1-031"  [ e:\�q�u���\1______________________�@�~\chapther2\031\sp031\031-schematic1-031.sim ] 

** Creating circuit file "031-schematic1-031.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\pwrmos.lib" 
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 101 0.1 10E9
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\031-SCHEMATIC1.net" 


.END
