** Profile: "SCHEMATIC1-s091_1"  [ C:\1________________________\chapther2\091\091-schematic1-s091_1.sim ] 

** Creating circuit file "091-schematic1-s091_1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "C:\Program Files\OrcadLite\Capture\Library\PSpice\siemens.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5.070U 0 0.5n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\091-SCHEMATIC1.net" 


.END
